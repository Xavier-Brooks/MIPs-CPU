library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use ieee.std_logic_unsigned.all;

entity Mem is
generic(mem_size : integer := 1024);
  Port (
        Addr :in std_logic_vector(27 downto 0);
        Dout :out std_logic_vector(31 downto 0)
        );
end Mem;

architecture beh of Mem is

Type MemT is array(0 to 2**17-1) of std_logic_vector(31 downto 0);
signal memory : MemT := (0 => "00100000000000010000000000000001", --puts the number 1 into R1
                         4 => "00100000000000100000000000000001", --puts 1 into R2
                         8 => "00100010000000000000000000000000", --NOP operation 
                         12 => "00100001111000000000000000000000",--NOP operation
                         16 => "00111100001000000000000000000001",--strs 1, 
                      --R1 + R2 = R3 
                         20 => "00000000001000100001100000100000",
                         24 => "00100010000000000000000000000000",--NOP operation 
                         28 => "00100001111000000000000000000000",--NOP operation
                         32 => "00111100010000000000000000000010",--strs 2
                      --R2 + R3 = R4
                         36 => "00000000010000110010000000100000",
                         40 => "00100010000000000000000000000000",--NOP operation 
                         44 => "00100001111000000000000000000000",--NOP operation
                         48 => "00111100011000000000000000000011",--strs 3
                      --R3 + R4 = R5    
                         52 => "00000000011001000010100000100000",
                         56 => "00100010000000000000000000000000",--NOP operation 
                         60 => "00100001111000000000000000000000",--NOP operation
                         64 => "00111100100000000000000000000101",--strs 5
                      --R4 + R5 = R6
                         68 => "00000000100001010011000000100000",
                         72 => "00100010000000000000000000000000",--NOP operation 
                         76 => "00100001111000000000000000000000",--NOP operation
                         80 => "00111100101000000000000000001000",--strs 8
                      --R5 + R6 = R7
                         84 => "00000000101001100011100000100000",
                         88 => "00100010000000000000000000000000",--NOP operation 
                         92 => "00100001111000000000000000000000",--NOP operation
                         96 => "00111100110000000000000000001101",--str 13
                      --R6 + R7 = R8
                         100 => "00000000110001110100000000100000",
                         104 => "00100010000000000000000000000000",--NOP operation 
                         108 => "00100001111000000000000000000000",--NOP operation
                         112 => "00111100111000000000000000010101",--str 21 
                      --R7 + R8 = R9
                         116 => "00000000111010000100100000100000",
                         120 => "00100010000000000000000000000000",--NOP operation 
                         124 => "00100001111000000000000000000000",--NOP operation
                         128 => "00111101000000000000000000100100",
                         
                      --R8 + R9 = R10    
                         132 => "00000001000010010101000000100000",
                         others => x"00000000");                      
begin 
     Dout <= memory(to_integer(unsigned(Addr(27 downto 0))));            
end beh;
